// top secret stuff
